-- +UEFSHDR----------------------------------------------------------------------
-- 2014 UEFS Universidade Estadual de Feira de Santana
-- TEC499-Sistemas Digitais
-- ------------------------------------------------------------------------------
-- TEAM: <Team identification>
-- ------------------------------------------------------------------------------
-- PROJECT: <Project Title>
-- ------------------------------------------------------------------------------
-- FILE NAME  : {module_name}
-- KEYWORDS 	: {keywords}
-- -----------------------------------------------------------------------------
-- PURPOSE: {description}
-- -UEFSHDR----------------------------------------------------------------------
